

module DE1_SoC_Computer (
	////////////////////////////////////
	// FPGA Pins
	////////////////////////////////////

	// Clock pins
	CLOCK_50,
	CLOCK2_50,
	CLOCK3_50,
	CLOCK4_50,

	// ADC
	ADC_CS_N,
	ADC_DIN,
	ADC_DOUT,
	ADC_SCLK,

	// Audio
	AUD_ADCDAT,
	AUD_ADCLRCK,
	AUD_BCLK,
	AUD_DACDAT,
	AUD_DACLRCK,
	AUD_XCK,

	// SDRAM
	DRAM_ADDR,
	DRAM_BA,
	DRAM_CAS_N,
	DRAM_CKE,
	DRAM_CLK,
	DRAM_CS_N,
	DRAM_DQ,
	DRAM_LDQM,
	DRAM_RAS_N,
	DRAM_UDQM,
	DRAM_WE_N,

	// I2C Bus for Configuration of the Audio and Video-In Chips
	FPGA_I2C_SCLK,
	FPGA_I2C_SDAT,

	// 40-Pin Headers
	GPIO_0,
	GPIO_1,
	
	// Seven Segment Displays
	HEX0,
	HEX1,
	HEX2,
	HEX3,
	HEX4,
	HEX5,

	// IR
	IRDA_RXD,
	IRDA_TXD,

	// Pushbuttons
	KEY,

	// LEDs
	LEDR,

	// PS2 Ports
	PS2_CLK,
	PS2_DAT,
	
	PS2_CLK2,
	PS2_DAT2,

	// Slider Switches
	SW,

	// Video-In
	TD_CLK27,
	TD_DATA,
	TD_HS,
	TD_RESET_N,
	TD_VS,

	// VGA
	VGA_B,
	VGA_BLANK_N,
	VGA_CLK,
	VGA_G,
	VGA_HS,
	VGA_R,
	VGA_SYNC_N,
	VGA_VS,

	////////////////////////////////////
	// HPS Pins
	////////////////////////////////////
	
	// DDR3 SDRAM
	HPS_DDR3_ADDR,
	HPS_DDR3_BA,
	HPS_DDR3_CAS_N,
	HPS_DDR3_CKE,
	HPS_DDR3_CK_N,
	HPS_DDR3_CK_P,
	HPS_DDR3_CS_N,
	HPS_DDR3_DM,
	HPS_DDR3_DQ,
	HPS_DDR3_DQS_N,
	HPS_DDR3_DQS_P,
	HPS_DDR3_ODT,
	HPS_DDR3_RAS_N,
	HPS_DDR3_RESET_N,
	HPS_DDR3_RZQ,
	HPS_DDR3_WE_N,

	// Ethernet
	HPS_ENET_GTX_CLK,
	HPS_ENET_INT_N,
	HPS_ENET_MDC,
	HPS_ENET_MDIO,
	HPS_ENET_RX_CLK,
	HPS_ENET_RX_DATA,
	HPS_ENET_RX_DV,
	HPS_ENET_TX_DATA,
	HPS_ENET_TX_EN,

	// Flash
	HPS_FLASH_DATA,
	HPS_FLASH_DCLK,
	HPS_FLASH_NCSO,

	// Accelerometer
	HPS_GSENSOR_INT,
		
	// General Purpose I/O
	HPS_GPIO,
		
	// I2C
	HPS_I2C_CONTROL,
	HPS_I2C1_SCLK,
	HPS_I2C1_SDAT,
	HPS_I2C2_SCLK,
	HPS_I2C2_SDAT,

	// Pushbutton
	HPS_KEY,

	// LED
	HPS_LED,
		
	// SD Card
	HPS_SD_CLK,
	HPS_SD_CMD,
	HPS_SD_DATA,

	// SPI
	HPS_SPIM_CLK,
	HPS_SPIM_MISO,
	HPS_SPIM_MOSI,
	HPS_SPIM_SS,

	// UART
	HPS_UART_RX,
	HPS_UART_TX,

	// USB
	HPS_CONV_USB_N,
	HPS_USB_CLKOUT,
	HPS_USB_DATA,
	HPS_USB_DIR,
	HPS_USB_NXT,
	HPS_USB_STP
);

//=======================================================
//  PARAMETER declarations
//=======================================================


//=======================================================
//  PORT declarations
//=======================================================

////////////////////////////////////
// FPGA Pins
////////////////////////////////////

// Clock pins
input						CLOCK_50;
input						CLOCK2_50;
input						CLOCK3_50;
input						CLOCK4_50;

// ADC
inout						ADC_CS_N;
output					ADC_DIN;
input						ADC_DOUT;
output					ADC_SCLK;

// Audio
input						AUD_ADCDAT;
inout						AUD_ADCLRCK;
inout						AUD_BCLK;
output					AUD_DACDAT;
inout						AUD_DACLRCK;
output					AUD_XCK;

// SDRAM
output 		[12: 0]	DRAM_ADDR;
output		[ 1: 0]	DRAM_BA;
output					DRAM_CAS_N;
output					DRAM_CKE;
output					DRAM_CLK;
output					DRAM_CS_N;
inout			[15: 0]	DRAM_DQ;
output					DRAM_LDQM;
output					DRAM_RAS_N;
output					DRAM_UDQM;
output					DRAM_WE_N;

// I2C Bus for Configuration of the Audio and Video-In Chips
output					FPGA_I2C_SCLK;
inout						FPGA_I2C_SDAT;

// 40-pin headers
inout			[35: 0]	GPIO_0;
inout			[35: 0]	GPIO_1;

// Seven Segment Displays
output		[ 6: 0]	HEX0;
output		[ 6: 0]	HEX1;
output		[ 6: 0]	HEX2;
output		[ 6: 0]	HEX3;
output		[ 6: 0]	HEX4;
output		[ 6: 0]	HEX5;

// IR
input						IRDA_RXD;
output					IRDA_TXD;

// Pushbuttons
input			[ 3: 0]	KEY;

// LEDs
output		[ 9: 0]	LEDR;

// PS2 Ports
inout						PS2_CLK;
inout						PS2_DAT;

inout						PS2_CLK2;
inout						PS2_DAT2;

// Slider Switches
input			[ 9: 0]	SW;

// Video-In
input						TD_CLK27;
input			[ 7: 0]	TD_DATA;
input						TD_HS;
output					TD_RESET_N;
input						TD_VS;

// VGA
output		[ 7: 0]	VGA_B;
output					VGA_BLANK_N;
output					VGA_CLK;
output		[ 7: 0]	VGA_G;
output					VGA_HS;
output		[ 7: 0]	VGA_R;
output					VGA_SYNC_N;
output					VGA_VS;



////////////////////////////////////
// HPS Pins
////////////////////////////////////
	
// DDR3 SDRAM
output		[14: 0]	HPS_DDR3_ADDR;
output		[ 2: 0]  HPS_DDR3_BA;
output					HPS_DDR3_CAS_N;
output					HPS_DDR3_CKE;
output					HPS_DDR3_CK_N;
output					HPS_DDR3_CK_P;
output					HPS_DDR3_CS_N;
output		[ 3: 0]	HPS_DDR3_DM;
inout			[31: 0]	HPS_DDR3_DQ;
inout			[ 3: 0]	HPS_DDR3_DQS_N;
inout			[ 3: 0]	HPS_DDR3_DQS_P;
output					HPS_DDR3_ODT;
output					HPS_DDR3_RAS_N;
output					HPS_DDR3_RESET_N;
input						HPS_DDR3_RZQ;
output					HPS_DDR3_WE_N;

// Ethernet
output					HPS_ENET_GTX_CLK;
inout						HPS_ENET_INT_N;
output					HPS_ENET_MDC;
inout						HPS_ENET_MDIO;
input						HPS_ENET_RX_CLK;
input			[ 3: 0]	HPS_ENET_RX_DATA;
input						HPS_ENET_RX_DV;
output		[ 3: 0]	HPS_ENET_TX_DATA;
output					HPS_ENET_TX_EN;

// Flash
inout			[ 3: 0]	HPS_FLASH_DATA;
output					HPS_FLASH_DCLK;
output					HPS_FLASH_NCSO;

// Accelerometer
inout						HPS_GSENSOR_INT;

// General Purpose I/O
inout			[ 1: 0]	HPS_GPIO;

// I2C
inout						HPS_I2C_CONTROL;
inout						HPS_I2C1_SCLK;
inout						HPS_I2C1_SDAT;
inout						HPS_I2C2_SCLK;
inout						HPS_I2C2_SDAT;

// Pushbutton
inout						HPS_KEY;

// LED
inout						HPS_LED;

// SD Card
output					HPS_SD_CLK;
inout						HPS_SD_CMD;
inout			[ 3: 0]	HPS_SD_DATA;

// SPI
output					HPS_SPIM_CLK;
input						HPS_SPIM_MISO;
output					HPS_SPIM_MOSI;
inout						HPS_SPIM_SS;

// UART
input						HPS_UART_RX;
output					HPS_UART_TX;

// USB
inout						HPS_CONV_USB_N;
input						HPS_USB_CLKOUT;
inout			[ 7: 0]	HPS_USB_DATA;
input						HPS_USB_DIR;
input						HPS_USB_NXT;
output					HPS_USB_STP;

//=======================================================
//  REG/WIRE declarations
//=======================================================

wire			[15: 0]	hex3_hex0;
//wire			[15: 0]	hex5_hex4;

//assign HEX0 = ~hex3_hex0[ 6: 0]; // hex3_hex0[ 6: 0]; 
//assign HEX1 = ~hex3_hex0[14: 8];
//assign HEX2 = ~hex3_hex0[22:16];
//assign HEX3 = ~hex3_hex0[30:24];
assign HEX4 = 7'b1111111;
assign HEX5 = 7'b1111111;

HexDigit Digit0(HEX0, hex3_hex0[3:0]);
HexDigit Digit1(HEX1, hex3_hex0[7:4]);
HexDigit Digit2(HEX2, hex3_hex0[11:8]);
HexDigit Digit3(HEX3, hex3_hex0[15:12]);

////=======================================================
//// Bus controller for AVALON bus-master
////=======================================================
//// computes DDS for sine wave and fills audio FIFO
//
//reg [31:0] bus_addr ; // Avalon address
//// see 
//// ftp://ftp.altera.com/up/pub/Altera_Material/15.1/University_Program_IP_Cores/Audio_Video/Audio.pdf
//// for addresses
//wire [31:0] audio_base_address = 32'h00003040 ;  // Avalon address
//wire [31:0] audio_fifo_address = 32'h00003044 ;  // Avalon address +4 offset
//wire [31:0] audio_left_address = 32'h00003048 ;  // Avalon address +8
//wire [31:0] audio_right_address = 32'h0000304c ;  // Avalon address +12
//reg [3:0] bus_byte_enable ; // four bit byte read/write mask
//reg bus_read  ;       // high when requesting data
//reg bus_write ;      //  high when writing data
//reg [31:0] bus_write_data ; //  data to send to Avalog bus
//wire bus_ack  ;       //  Avalon bus raises this when done
//wire [31:0] bus_read_data ; // data from Avalon bus
//reg [30:0] timer ;
//reg [3:0] state ;
//wire state_clock ;
//
//// current free words in audio interface
//reg [7:0] fifo_space ;
//// debug check of space
//assign LEDR = fifo_space ;
//
//// use 4-byte-wide bus-master	 
////assign bus_byte_enable = 4'b1111;
//
//// DDS signals
//reg [31:0] dds_accum ;
//// DDS LUT
//wire [15:0] sine_out ;
//sync_rom sineTable(CLOCK_50, dds_accum[31:24], sine_out);
//
//// get some signals exposed
//// connect bus master signals to i/o for probes
//assign GPIO_0[0] = bus_write ;
//assign GPIO_0[1] = bus_read ;
//assign GPIO_0[2] = bus_ack ;
////assign GPIO_0[3] = ??? ;
//
//
//
//always @(posedge CLOCK_50) begin //CLOCK_50
//
//	// reset state machine and read/write controls
//	if (~KEY[0]) begin
//		state <= 0 ;
//		bus_read <= 0 ; // set to one if a read opeation from bus
//		bus_write <= 0 ; // set to one if a write operation to bus
//		timer <= 0;
//	end
//	else begin
//		// timer just for deubgging
//		timer <= timer + 1;
//	end
//	
//	// set up read FIFO available space
//	if (state==4'd0) begin
//		bus_addr <= audio_fifo_address ;
//		bus_read <= 1'b1 ;
//		bus_byte_enable <= 4'b1111;
//		state <= 4'd1 ; // wait for read ACK
//	end
//	
//	// wait for read ACK and read the fifo available
//	// bus ACK is high when data is available
//	if (state==4'd1 && bus_ack==1) begin
//		state <= 4'd2 ; //4'd2
//		// FIFO space is in high byte
//		fifo_space <= (bus_read_data>>24) ;
//		// end the read
//		bus_read <= 1'b0 ;
//	end
//	
//	// When there is room in the FIFO
//	// -- compute next DDS sine sample
//	// -- start write to fifo for each channel
//	// -- first the left channel
//	if (state==4'd2 && fifo_space>8'd2) begin // 
//		state <= 4'd3;	
//		// IF SW=10'h200 
//		// and Fout = (sample_rate)/(2^32)*{SW[9:0], 16'b0}
//		// then Fout=48000/(2^32)*(2^25) = 375 Hz
//		dds_accum <= dds_accum + {SW[9:0], 16'b0} ;
//		// convert 16-bit table to 32-bit format
//		bus_write_data <= (sine_out << 16) ;
//		bus_addr <= audio_left_address ;
//		bus_byte_enable <= 4'b1111;
//		bus_write <= 1'b1 ;
//	end	
//	// if no space, try again later
//	else if (state==4'd2 && fifo_space<=8'd2) begin
//		state <= 4'b0 ;
//	end
//	
//	// detect bus-transaction-complete ACK 
//	// for left channel write
//	// You MUST do this check
//	if (state==4'd3 && bus_ack==1) begin
//		state <= 4'd4 ;
//		bus_write <= 0;
//	end
//	
//	// -- now the right channel
//	if (state==4'd4) begin // 
//		state <= 4'd5;	
//		bus_write_data <= (sine_out << 16) ;
//		bus_addr <= audio_right_address ;
//		bus_write <= 1'b1 ;
//	end	
//	
//	// detect bus-transaction-complete ACK
//	// for right channel write
//	// You MUST do this check
//	if (state==4'd5 && bus_ack==1) begin
//		state <= 4'd0 ;
//		bus_write <= 0;
//	end
//	
//end // always @(posedge state_clock)


//=======================================================
// Integrator DDS
//=======================================================


// see 
// ftp://ftp.altera.com/up/pub/Altera_Material/15.1/University_Program_IP_Cores/Audio_Video/Audio.pdf
// for addresses
wire [31:0] audio_base_address = 32'h00003040 ;  // Avalon address
wire [31:0] audio_fifo_address = 32'h00003044 ;  // Avalon address +4 offset
wire [31:0] audio_left_address = 32'h00003048 ;  // Avalon address +8
wire [31:0] audio_right_address = 32'h0000304c ;  // Avalon address +12

wire state_clock ;


// use 4-byte-wide bus-master	 
//assign bus_byte_enable = 4'b1111;

// get some signals exposed
// connect bus master signals to i/o for probes
assign GPIO_0[0] = bus_write ;
assign GPIO_0[1] = bus_read ;
assign GPIO_0[2] = bus_ack ;
//assign GPIO_0[3] = ??? ;

reg [3:0] state ;
reg bus_read  ;       // high when requesting data
reg bus_write ;      //  high when writing data
reg [30:0] timer ;

reg [31:0] bus_addr ; // Avalon address
reg [3:0] bus_byte_enable ; // four bit byte read/write mask

wire bus_ack  ;       //  Avalon bus raises this when done
wire [31:0] bus_read_data ; // data from Avalon bus

// current free words in audio interface
reg [7:0] fifo_space ;


// debug check of space
assign LEDR = fifo_space ;


reg [31:0] bus_write_data ; //  data to send to Avalog bus

// DDS signals
reg [31:0] dds_accum_x, dds_accum_y, dds_accum_z;

wire [31:0] dds_incr_x, dds_incr_y, dds_incr_z;

wire [15:0] sine_out_x, sine_out_y, sine_out_z;

wire [31:0] sine_ext_x, sine_ext_y, sine_ext_z;

assign sine_ext_x = { {16{sine_out_x[15]}}, sine_out_x };
assign sine_ext_y = { {16{sine_out_y[15]}}, sine_out_y };
assign sine_ext_z = { {16{sine_out_z[15]}}, sine_out_z };

freq_LUT DDS_x (
	.address( testbench_out_x[25:20] ),
	.dds_increment_out( dds_incr_x )
);

freq_LUT DDS_y (
	.address( testbench_out_y[25:20] ),
	.dds_increment_out( dds_incr_y )
);

freq_LUT DDS_z (
	.address( testbench_out_z[25:20] ),
	.dds_increment_out( dds_incr_z )
);

sync_rom sine_x (
	.clock(CLOCK_50), 
	.address(dds_accum_x[31:24]), 
	.sine(sine_out_x)
);

sync_rom sine_y (
	.clock(CLOCK_50), 
	.address(dds_accum_y[31:24]), 
	.sine(sine_out_y)
);

sync_rom sine_z (
	.clock(CLOCK_50), 
	.address(dds_accum_z[31:24]), 
	.sine(sine_out_z)
);


always @(posedge CLOCK_50) begin //CLOCK_50

	// reset state machine and read/write controls
	if (arm_reset[0] == 0) begin
		state <= 0 ;
		bus_read <= 0 ; // set to one if a read opeation from bus
		bus_write <= 0 ; // set to one if a write operation to bus
		timer <= 0;
	end
	else begin
		// timer just for deubgging
		timer <= timer + 1;
	end
	
	// set up read FIFO available space
	if (state==4'd0) begin
		bus_addr <= audio_fifo_address ;
		bus_read <= 1'b1 ;
		bus_byte_enable <= 4'b1111;
		state <= 4'd1 ; // wait for read ACK
	end
	
	// wait for read ACK and read the fifo available
	// bus ACK is high when data is available
	if (state==4'd1 && bus_ack==1) begin
		state <= 4'd2 ; //4'd2
		// FIFO space is in high byte
		fifo_space <= (bus_read_data>>24) ;
		// end the read
		bus_read <= 1'b0 ;
	end
	
	// When there is room in the FIFO
	// -- compute next DDS sine sample
	// -- start write to fifo for each channel
	// -- first the left channel
	if (state==4'd2 && fifo_space>8'd2) begin // 
		state <= 4'd3;	
		// IF SW=10'h200 
		// and Fout = (sample_rate)/(2^32)*{SW[9:0], 16'b0}
		// then Fout=48000/(2^32)*(2^25) = 375 Hz
		dds_accum_x <= dds_accum_x + dds_incr_x ;
		dds_accum_y <= dds_accum_y + dds_incr_y ;
		dds_accum_z <= dds_accum_z + dds_incr_z ;
		// convert 16-bit table to 32-bit format
		bus_write_data <= (sine_ext_x << 14) + (sine_ext_y << 14) + (sine_ext_z << 14);
		bus_addr <= audio_left_address ;
		bus_byte_enable <= 4'b1111;
		bus_write <= 1'b1 ;
	end	
	// if no space, try again later
	else if (state==4'd2 && fifo_space<=8'd2) begin
		state <= 4'b0 ;
	end
	
	// detect bus-transaction-complete ACK 
	// for left channel write
	// You MUST do this check
	if (state==4'd3 && bus_ack==1) begin
		state <= 4'd4 ;
		bus_write <= 0;
	end
	
	// -- now the right channel
	if (state==4'd4) begin // 
		state <= 4'd5;	
		bus_write_data <= (sine_ext_x << 14) + (sine_ext_y << 14) + (sine_ext_z << 14);
		bus_addr <= audio_right_address ;
		bus_write <= 1'b1 ;
	end	
	
	// detect bus-transaction-complete ACK
	// for right channel write
	// You MUST do this check
	if (state==4'd5 && bus_ack==1) begin
		state <= 4'd0 ;
		bus_write <= 0;
	end
	
end // always @(posedge state_clock)


//=======================================================
// DDA Stuff
//=======================================================


wire signed [26:0] testbench_out_x, testbench_out_y, testbench_out_z;
wire signed [31:0] dt_val, x_val, y_val, z_val, sig_val, beta_val, rho_val;
wire signed [31:0] signed_x, signed_y, signed_z;
wire [7:0]         arm_clock, arm_reset, start_stop;

DDA DUT (
	  .clock(arm_clock[0]), 
	  .reset(arm_reset[0]), 
	  .dt_init( { 27'b0000000_00000001000000000000 } ),
	  .x_init( x_val[26:0] ),
	  .y_init( y_val[26:0] ),
	  .z_init( z_val[26:0] ),
	  .sigma_init( sig_val[26:0] ),
	  .rho_init( rho_val[26:0] ),
	  .beta_init( beta_val[26:0] ),
	  .out_x(testbench_out_x),
	  .out_y(testbench_out_y),
	  .out_z(testbench_out_z),
	  .start_stop(start_stop[0])
);

assign signed_x = { {5{testbench_out_x[26]}}, testbench_out_x };
assign signed_y = { {5{testbench_out_y[26]}}, testbench_out_y };
assign signed_z = { {5{testbench_out_z[26]}}, testbench_out_z };

//=======================================================
//  Structural coding
//=======================================================

Computer_System The_System (
	////////////////////////////////////
	// FPGA Side
	////////////////////////////////////

	// Global signals
	.system_pll_ref_clk_clk					(CLOCK_50),
	.system_pll_ref_reset_reset			(1'b0),

	// AV Config
	.av_config_SCLK							(FPGA_I2C_SCLK),
	.av_config_SDAT							(FPGA_I2C_SDAT),
	
	// Audio Subsystem
	.audio_pll_ref_clk_clk					(CLOCK3_50),
	.audio_pll_ref_reset_reset				(1'b0),
	.audio_clk_clk								(AUD_XCK),
	.audio_ADCDAT								(AUD_ADCDAT),
	.audio_ADCLRCK								(AUD_ADCLRCK),
	.audio_BCLK									(AUD_BCLK),
	.audio_DACDAT								(AUD_DACDAT),
	.audio_DACLRCK								(AUD_DACLRCK),
	
	// bus-master state machine interface
	.bus_master_audio_external_interface_address     (bus_addr),     
	.bus_master_audio_external_interface_byte_enable (bus_byte_enable), 
	.bus_master_audio_external_interface_read        (bus_read),        
	.bus_master_audio_external_interface_write       (bus_write),       
	.bus_master_audio_external_interface_write_data  (bus_write_data),  
	.bus_master_audio_external_interface_acknowledge (bus_ack),                                  
	.bus_master_audio_external_interface_read_data   (bus_read_data),  

	// VGA Subsystem
	.vga_pll_ref_clk_clk 					(CLOCK2_50),
	.vga_pll_ref_reset_reset				(1'b0),
	.vga_CLK										(VGA_CLK),
	.vga_BLANK									(VGA_BLANK_N),
	.vga_SYNC									(VGA_SYNC_N),
	.vga_HS										(VGA_HS),
	.vga_VS										(VGA_VS),
	.vga_R										(VGA_R),
	.vga_G										(VGA_G),
	.vga_B										(VGA_B),
	
	// SDRAM
	.sdram_clk_clk								(DRAM_CLK),
   .sdram_addr									(DRAM_ADDR),
	.sdram_ba									(DRAM_BA),
	.sdram_cas_n								(DRAM_CAS_N),
	.sdram_cke									(DRAM_CKE),
	.sdram_cs_n									(DRAM_CS_N),
	.sdram_dq									(DRAM_DQ),
	.sdram_dqm									({DRAM_UDQM,DRAM_LDQM}),
	.sdram_ras_n								(DRAM_RAS_N),
	.sdram_we_n									(DRAM_WE_N),
	
	// Solver Subsystem
	.x_pio_ext_export                   (signed_x),
	.y_pio_ext_export                   (signed_y),
	.z_pio_ext_export                   (signed_z),
   .plot_clock_ext_export              (arm_clock),
	.plot_reset_ext_export              (arm_reset),
	.x_init_pio_ext_export              (x_val),
	.y_init_pio_ext_export              (y_val),
	.z_init_pio_ext_export              (z_val),
	.sig_pio_ext_export                 (sig_val),
	.rho_pio_ext_export                 (rho_val),
	.beta_pio_ext_export                (beta_val),
	.start_stop_pio_ext_export          (start_stop),
	
	////////////////////////////////////
	// HPS Side
	////////////////////////////////////
	// DDR3 SDRAM
	.memory_mem_a			(HPS_DDR3_ADDR),
	.memory_mem_ba			(HPS_DDR3_BA),
	.memory_mem_ck			(HPS_DDR3_CK_P),
	.memory_mem_ck_n		(HPS_DDR3_CK_N),
	.memory_mem_cke		(HPS_DDR3_CKE),
	.memory_mem_cs_n		(HPS_DDR3_CS_N),
	.memory_mem_ras_n		(HPS_DDR3_RAS_N),
	.memory_mem_cas_n		(HPS_DDR3_CAS_N),
	.memory_mem_we_n		(HPS_DDR3_WE_N),
	.memory_mem_reset_n	(HPS_DDR3_RESET_N),
	.memory_mem_dq			(HPS_DDR3_DQ),
	.memory_mem_dqs		(HPS_DDR3_DQS_P),
	.memory_mem_dqs_n		(HPS_DDR3_DQS_N),
	.memory_mem_odt		(HPS_DDR3_ODT),
	.memory_mem_dm			(HPS_DDR3_DM),
	.memory_oct_rzqin		(HPS_DDR3_RZQ),
		  
	// Ethernet
	.hps_io_hps_io_gpio_inst_GPIO35	(HPS_ENET_INT_N),
	.hps_io_hps_io_emac1_inst_TX_CLK	(HPS_ENET_GTX_CLK),
	.hps_io_hps_io_emac1_inst_TXD0	(HPS_ENET_TX_DATA[0]),
	.hps_io_hps_io_emac1_inst_TXD1	(HPS_ENET_TX_DATA[1]),
	.hps_io_hps_io_emac1_inst_TXD2	(HPS_ENET_TX_DATA[2]),
	.hps_io_hps_io_emac1_inst_TXD3	(HPS_ENET_TX_DATA[3]),
	.hps_io_hps_io_emac1_inst_RXD0	(HPS_ENET_RX_DATA[0]),
	.hps_io_hps_io_emac1_inst_MDIO	(HPS_ENET_MDIO),
	.hps_io_hps_io_emac1_inst_MDC		(HPS_ENET_MDC),
	.hps_io_hps_io_emac1_inst_RX_CTL	(HPS_ENET_RX_DV),
	.hps_io_hps_io_emac1_inst_TX_CTL	(HPS_ENET_TX_EN),
	.hps_io_hps_io_emac1_inst_RX_CLK	(HPS_ENET_RX_CLK),
	.hps_io_hps_io_emac1_inst_RXD1	(HPS_ENET_RX_DATA[1]),
	.hps_io_hps_io_emac1_inst_RXD2	(HPS_ENET_RX_DATA[2]),
	.hps_io_hps_io_emac1_inst_RXD3	(HPS_ENET_RX_DATA[3]),

	// Flash
	.hps_io_hps_io_qspi_inst_IO0	(HPS_FLASH_DATA[0]),
	.hps_io_hps_io_qspi_inst_IO1	(HPS_FLASH_DATA[1]),
	.hps_io_hps_io_qspi_inst_IO2	(HPS_FLASH_DATA[2]),
	.hps_io_hps_io_qspi_inst_IO3	(HPS_FLASH_DATA[3]),
	.hps_io_hps_io_qspi_inst_SS0	(HPS_FLASH_NCSO),
	.hps_io_hps_io_qspi_inst_CLK	(HPS_FLASH_DCLK),

	// Accelerometer
	.hps_io_hps_io_gpio_inst_GPIO61	(HPS_GSENSOR_INT),

	//.adc_sclk                        (ADC_SCLK),
	//.adc_cs_n                        (ADC_CS_N),
	//.adc_dout                        (ADC_DOUT),
	//.adc_din                         (ADC_DIN),

	// General Purpose I/O
	.hps_io_hps_io_gpio_inst_GPIO40	(HPS_GPIO[0]),
	.hps_io_hps_io_gpio_inst_GPIO41	(HPS_GPIO[1]),

	// I2C
	.hps_io_hps_io_gpio_inst_GPIO48	(HPS_I2C_CONTROL),
	.hps_io_hps_io_i2c0_inst_SDA		(HPS_I2C1_SDAT),
	.hps_io_hps_io_i2c0_inst_SCL		(HPS_I2C1_SCLK),
	.hps_io_hps_io_i2c1_inst_SDA		(HPS_I2C2_SDAT),
	.hps_io_hps_io_i2c1_inst_SCL		(HPS_I2C2_SCLK),

	// Pushbutton
	.hps_io_hps_io_gpio_inst_GPIO54	(HPS_KEY),

	// LED
	.hps_io_hps_io_gpio_inst_GPIO53	(HPS_LED),

	// SD Card
	.hps_io_hps_io_sdio_inst_CMD	(HPS_SD_CMD),
	.hps_io_hps_io_sdio_inst_D0	(HPS_SD_DATA[0]),
	.hps_io_hps_io_sdio_inst_D1	(HPS_SD_DATA[1]),
	.hps_io_hps_io_sdio_inst_CLK	(HPS_SD_CLK),
	.hps_io_hps_io_sdio_inst_D2	(HPS_SD_DATA[2]),
	.hps_io_hps_io_sdio_inst_D3	(HPS_SD_DATA[3]),

	// SPI
	.hps_io_hps_io_spim1_inst_CLK		(HPS_SPIM_CLK),
	.hps_io_hps_io_spim1_inst_MOSI	(HPS_SPIM_MOSI),
	.hps_io_hps_io_spim1_inst_MISO	(HPS_SPIM_MISO),
	.hps_io_hps_io_spim1_inst_SS0		(HPS_SPIM_SS),

	// UART
	.hps_io_hps_io_uart0_inst_RX	(HPS_UART_RX),
	.hps_io_hps_io_uart0_inst_TX	(HPS_UART_TX),

	// USB
	.hps_io_hps_io_gpio_inst_GPIO09	(HPS_CONV_USB_N),
	.hps_io_hps_io_usb1_inst_D0		(HPS_USB_DATA[0]),
	.hps_io_hps_io_usb1_inst_D1		(HPS_USB_DATA[1]),
	.hps_io_hps_io_usb1_inst_D2		(HPS_USB_DATA[2]),
	.hps_io_hps_io_usb1_inst_D3		(HPS_USB_DATA[3]),
	.hps_io_hps_io_usb1_inst_D4		(HPS_USB_DATA[4]),
	.hps_io_hps_io_usb1_inst_D5		(HPS_USB_DATA[5]),
	.hps_io_hps_io_usb1_inst_D6		(HPS_USB_DATA[6]),
	.hps_io_hps_io_usb1_inst_D7		(HPS_USB_DATA[7]),
	.hps_io_hps_io_usb1_inst_CLK		(HPS_USB_CLKOUT),
	.hps_io_hps_io_usb1_inst_STP		(HPS_USB_STP),
	.hps_io_hps_io_usb1_inst_DIR		(HPS_USB_DIR),
	.hps_io_hps_io_usb1_inst_NXT		(HPS_USB_NXT)
);


endmodule

/////////////////////////////////////////////////
//// DDA ////////////////////////////////////////
/////////////////////////////////////////////////

module DDA (
    clock, 
    reset, 
    dt_init, 
    x_init, 
    y_init, 
    z_init,
    sigma_init,
    rho_init,
    beta_init,
    out_x,
    out_y,
    out_z,
	 start_stop );

    input  signed clock, reset, start_stop;
    input  signed [26:0] dt_init, x_init, y_init, z_init, sigma_init, rho_init, beta_init;
    output signed [26:0] out_x, out_y, out_z;

    wire signed [26:0] int_out_x, int_out_y, int_out_z, dxdt_out, dydt_out, dzdt_out;

    dxdt dxdt_inst (
        .out(dxdt_out), 
        .sigma(sigma_init),
        .x_(int_out_x),
        .y_(int_out_y),
        .dt(dt_init)
    );

    dydt dydt_inst (
        .out(dydt_out), 
        .rho(rho_init),
        .x_(int_out_x),
        .y_(int_out_y),
        .z_(int_out_z),
        .dt(dt_init)
    );

    dzdt dzdt_inst (
        .out(dzdt_out), 
        .beta(beta_init),
        .x_(int_out_x),
        .y_(int_out_y),
        .z_(int_out_z),
        .dt(dt_init)
    );

    integrator int_inst_x (
        .out(int_out_x), 
        .funct(dxdt_out), 
        .InitialOut(x_init),
        .clk(clock),
        .reset(reset),
		  .start_stop(start_stop)
    );

    integrator int_inst_y (
        .out(int_out_y), 
        .funct(dydt_out), 
        .InitialOut(y_init),
        .clk(clock),
        .reset(reset),
		  .start_stop(start_stop)
    );

    integrator int_inst_z (
        .out(int_out_z), 
        .funct(dzdt_out), 
        .InitialOut(z_init),
        .clk(clock),
        .reset(reset),
		  .start_stop(start_stop)
    );

    assign out_x = int_out_x;
    assign out_y = int_out_y;
    assign out_z = int_out_z;

endmodule

/////////////////////////////////////////////////
//// funct: dx*dt ///////////////////////////////
/////////////////////////////////////////////////

module dxdt (out, sigma, x_, y_, dt);
	output signed [26:0] out;  // fed into integrator
	input  signed [26:0] sigma;
	input  signed [26:0] x_, y_, dt;
	
	wire signed	  [26:0] mult_out1, dt_mult, y_sub_x;

    assign y_sub_x = y_ - x_;
    assign dt_mult = y_sub_x >>> 8;
	signed_mult sign_mult_sigma (.out(mult_out1), .a(sigma), .b(dt_mult));
    assign out = mult_out1;

endmodule

/////////////////////////////////////////////////
//// funct: dy*dt ///////////////////////////////
/////////////////////////////////////////////////

module dydt (out, rho, x_, y_, z_, dt);
	output signed [26:0] out;  // fed into integrator
	input  signed [26:0] rho;
	input  signed [26:0] x_, y_, z_, dt;
	
	wire signed	  [26:0] mult_out1, rho_sub_z, dt_mult_rho_z, dt_mult_y;

    assign rho_sub_z = rho - z_;
    assign dt_mult_rho_z = rho_sub_z >>> 8;
    assign dt_mult_y = y_ >>> 8;
	signed_mult sign_mult_x (.out(mult_out1), .a(x_), .b(dt_mult_rho_z));
    assign out = mult_out1 - dt_mult_y;

endmodule

/////////////////////////////////////////////////
//// funct: dz*dt ///////////////////////////////
/////////////////////////////////////////////////

module dzdt (out, beta, x_, y_, z_, dt);
	output signed [26:0] out;  // fed into integrator
	input  signed [26:0] beta;
	input  signed [26:0] x_, y_, z_, dt;
	
	wire signed	  [26:0] mult_x_y, mult_beta_z, dt_mult_y, dt_mult_z;

    assign dt_mult_y = y_ >>> 8;
    assign dt_mult_z = z_ >>> 8;

	signed_mult sign_mult_x_y (.out(mult_x_y), .a(x_), .b(dt_mult_y));
    signed_mult sign_mult_beta_z (.out(mult_beta_z), .a(beta), .b(dt_mult_z));
    assign out = mult_x_y - mult_beta_z;

endmodule

/////////////////////////////////////////////////
//// general integrator /////////////////////////
/////////////////////////////////////////////////

module integrator (out, funct, InitialOut, clk, reset, start_stop);
	output signed [26:0] out; 		 // the state variable V
	input  signed [26:0] funct;      // the dV/dt function
	input  clk, reset, start_stop;
	input  signed [26:0] InitialOut;  // the initial state variable V
	
	wire signed	[26:0] out, v1new;
	reg  signed	[26:0] v1;
	
	always @ (posedge clk) begin
		if (reset == 0)
			v1 <= InitialOut;
		else if (start_stop == 0)
			v1 <= v1new;	
		else
			v1 <= v1;
	end

	assign v1new = v1 + funct;
	assign out = v1;

endmodule

//////////////////////////////////////////////////
//// signed mult of 7.20 format 2'comp////////////
//////////////////////////////////////////////////

module signed_mult (out, a, b);
	output 	signed  [26:0]	out;
	input 	signed	[26:0] 	a;
	input 	signed	[26:0] 	b;
	// intermediate full bit length
	wire 	signed	[53:0]	mult_out;
	assign mult_out = a * b;
	// select bits for 7.20 fixed point
	assign out = { mult_out[53], mult_out[45:20] };

endmodule

//////////////////////////////////////////////////

//////////////////////////////////////////////////
////////////	DDS FOR INTEGRATOR	//////////////
//////////////////////////////////////////////////

module freq_LUT (
    input wire [5:0] address,
    output wire [31:0] dds_increment_out
);
reg [31:0] dds_increment ; 
always@(address)
begin
    case(address)
        6'd0: dds_increment=32'd2460658;
        6'd1: dds_increment=32'd2762200;
        6'd2: dds_increment=32'd2925946;
        6'd3: dds_increment=32'd3284755;
        6'd4: dds_increment=32'd3686513;
        6'd5: dds_increment=32'd3905735;
        6'd6: dds_increment=32'd4384445;
        6'd7: dds_increment=32'd4921316;
        6'd8: dds_increment=32'd5524401;
        6'd9: dds_increment=32'd5852787;
        6'd10: dds_increment=32'd6569510;
        6'd11: dds_increment=32'd7373921;
        6'd12: dds_increment=32'd7812366;
        6'd13: dds_increment=32'd8768891;
        6'd14: dds_increment=32'd9842633;
        6'd15: dds_increment=32'd11047908;
        6'd16: dds_increment=32'd11704680;
        6'd17: dds_increment=32'd13138126;
        6'd18: dds_increment=32'd14746949;
        6'd19: dds_increment=32'd15623838;
        6'd20: dds_increment=32'd17537783;
        6'd21: dds_increment=32'd19685266;
        6'd22: dds_increment=32'd22095817;
        6'd23: dds_increment=32'd23410256;
        6'd24: dds_increment=32'd26276252;
        6'd25: dds_increment=32'd29494793;
        6'd26: dds_increment=32'd31248571;
        6'd27: dds_increment=32'd35075566;
        6'd28: dds_increment=32'd39370533;
        6'd29: dds_increment=32'd44191634;
        6'd30: dds_increment=32'd46819617;
        6'd31: dds_increment=32'd52553398;
        6'd32: dds_increment=32'd58988691;
        6'd33: dds_increment=32'd62497142;
        6'd34: dds_increment=32'd70150237;
        6'd35: dds_increment=32'd78741067;
        6'd36: dds_increment=32'd88384163;
        6'd37: dds_increment=32'd93639234;
        6'd38: dds_increment=32'd105106797;
        6'd39: dds_increment=32'd117978277;
        6'd40: dds_increment=32'd124993390;
        6'd41: dds_increment=32'd140300475;
        6'd42: dds_increment=32'd157482134;
        6'd43: dds_increment=32'd176767432;
        6'd44: dds_increment=32'd187278469;
        6'd45: dds_increment=32'd210213595;
        6'd46: dds_increment=32'd235956555;
        6'd47: dds_increment=32'd249987676;
        6'd48: dds_increment=32'd280600950;
        6'd49: dds_increment=32'd314964268;
        6'd50: dds_increment=32'd353535759;
        6'd51: dds_increment=32'd374557834;
        default dds_increment =32'd0 ;
    endcase
end
assign dds_increment_out = dds_increment ;
endmodule


//////////////////////////////////////////////////
////////////	Sin Wave ROM Table	//////////////
//////////////////////////////////////////////////
// produces a 2's comp, 16-bit, approximation
// of a sine wave, given an input phase (address)
module sync_rom (clock, address, sine);
input clock;
input [7:0] address;
output [15:0] sine;
reg signed [15:0] sine;
always@(posedge clock)
begin
    case(address)
    		8'h00: sine = 16'h0000 ;
			8'h01: sine = 16'h0192 ;
			8'h02: sine = 16'h0323 ;
			8'h03: sine = 16'h04b5 ;
			8'h04: sine = 16'h0645 ;
			8'h05: sine = 16'h07d5 ;
			8'h06: sine = 16'h0963 ;
			8'h07: sine = 16'h0af0 ;
			8'h08: sine = 16'h0c7c ;
			8'h09: sine = 16'h0e05 ;
			8'h0a: sine = 16'h0f8c ;
			8'h0b: sine = 16'h1111 ;
			8'h0c: sine = 16'h1293 ;
			8'h0d: sine = 16'h1413 ;
			8'h0e: sine = 16'h158f ;
			8'h0f: sine = 16'h1708 ;
			8'h10: sine = 16'h187d ;
			8'h11: sine = 16'h19ef ;
			8'h12: sine = 16'h1b5c ;
			8'h13: sine = 16'h1cc5 ;
			8'h14: sine = 16'h1e2a ;
			8'h15: sine = 16'h1f8b ;
			8'h16: sine = 16'h20e6 ;
			8'h17: sine = 16'h223c ;
			8'h18: sine = 16'h238d ;
			8'h19: sine = 16'h24d9 ;
			8'h1a: sine = 16'h261f ;
			8'h1b: sine = 16'h275f ;
			8'h1c: sine = 16'h2899 ;
			8'h1d: sine = 16'h29cc ;
			8'h1e: sine = 16'h2afa ;
			8'h1f: sine = 16'h2c20 ;
			8'h20: sine = 16'h2d40 ;
			8'h21: sine = 16'h2e59 ;
			8'h22: sine = 16'h2f6b ;
			8'h23: sine = 16'h3075 ;
			8'h24: sine = 16'h3178 ;
			8'h25: sine = 16'h3273 ;
			8'h26: sine = 16'h3366 ;
			8'h27: sine = 16'h3452 ;
			8'h28: sine = 16'h3535 ;
			8'h29: sine = 16'h3611 ;
			8'h2a: sine = 16'h36e4 ;
			8'h2b: sine = 16'h37ae ;
			8'h2c: sine = 16'h3870 ;
			8'h2d: sine = 16'h3929 ;
			8'h2e: sine = 16'h39da ;
			8'h2f: sine = 16'h3a81 ;
			8'h30: sine = 16'h3b1f ;
			8'h31: sine = 16'h3bb5 ;
			8'h32: sine = 16'h3c41 ;
			8'h33: sine = 16'h3cc4 ;
			8'h34: sine = 16'h3d3d ;
			8'h35: sine = 16'h3dad ;
			8'h36: sine = 16'h3e14 ;
			8'h37: sine = 16'h3e70 ;
			8'h38: sine = 16'h3ec4 ;
			8'h39: sine = 16'h3f0d ;
			8'h3a: sine = 16'h3f4d ;
			8'h3b: sine = 16'h3f83 ;
			8'h3c: sine = 16'h3fb0 ;
			8'h3d: sine = 16'h3fd2 ;
			8'h3e: sine = 16'h3feb ;
			8'h3f: sine = 16'h3ffa ;
			8'h40: sine = 16'h3fff ;
			8'h41: sine = 16'h3ffa ;
			8'h42: sine = 16'h3feb ;
			8'h43: sine = 16'h3fd2 ;
			8'h44: sine = 16'h3fb0 ;
			8'h45: sine = 16'h3f83 ;
			8'h46: sine = 16'h3f4d ;
			8'h47: sine = 16'h3f0d ;
			8'h48: sine = 16'h3ec4 ;
			8'h49: sine = 16'h3e70 ;
			8'h4a: sine = 16'h3e14 ;
			8'h4b: sine = 16'h3dad ;
			8'h4c: sine = 16'h3d3d ;
			8'h4d: sine = 16'h3cc4 ;
			8'h4e: sine = 16'h3c41 ;
			8'h4f: sine = 16'h3bb5 ;
			8'h50: sine = 16'h3b1f ;
			8'h51: sine = 16'h3a81 ;
			8'h52: sine = 16'h39da ;
			8'h53: sine = 16'h3929 ;
			8'h54: sine = 16'h3870 ;
			8'h55: sine = 16'h37ae ;
			8'h56: sine = 16'h36e4 ;
			8'h57: sine = 16'h3611 ;
			8'h58: sine = 16'h3535 ;
			8'h59: sine = 16'h3452 ;
			8'h5a: sine = 16'h3366 ;
			8'h5b: sine = 16'h3273 ;
			8'h5c: sine = 16'h3178 ;
			8'h5d: sine = 16'h3075 ;
			8'h5e: sine = 16'h2f6b ;
			8'h5f: sine = 16'h2e59 ;
			8'h60: sine = 16'h2d40 ;
			8'h61: sine = 16'h2c20 ;
			8'h62: sine = 16'h2afa ;
			8'h63: sine = 16'h29cc ;
			8'h64: sine = 16'h2899 ;
			8'h65: sine = 16'h275f ;
			8'h66: sine = 16'h261f ;
			8'h67: sine = 16'h24d9 ;
			8'h68: sine = 16'h238d ;
			8'h69: sine = 16'h223c ;
			8'h6a: sine = 16'h20e6 ;
			8'h6b: sine = 16'h1f8b ;
			8'h6c: sine = 16'h1e2a ;
			8'h6d: sine = 16'h1cc5 ;
			8'h6e: sine = 16'h1b5c ;
			8'h6f: sine = 16'h19ef ;
			8'h70: sine = 16'h187d ;
			8'h71: sine = 16'h1708 ;
			8'h72: sine = 16'h158f ;
			8'h73: sine = 16'h1413 ;
			8'h74: sine = 16'h1293 ;
			8'h75: sine = 16'h1111 ;
			8'h76: sine = 16'h0f8c ;
			8'h77: sine = 16'h0e05 ;
			8'h78: sine = 16'h0c7c ;
			8'h79: sine = 16'h0af0 ;
			8'h7a: sine = 16'h0963 ;
			8'h7b: sine = 16'h07d5 ;
			8'h7c: sine = 16'h0645 ;
			8'h7d: sine = 16'h04b5 ;
			8'h7e: sine = 16'h0323 ;
			8'h7f: sine = 16'h0192 ;
			8'h80: sine = 16'h0000 ;
			8'h81: sine = 16'hfe6e ;
			8'h82: sine = 16'hfcdd ;
			8'h83: sine = 16'hfb4b ;
			8'h84: sine = 16'hf9bb ;
			8'h85: sine = 16'hf82b ;
			8'h86: sine = 16'hf69d ;
			8'h87: sine = 16'hf510 ;
			8'h88: sine = 16'hf384 ;
			8'h89: sine = 16'hf1fb ;
			8'h8a: sine = 16'hf074 ;
			8'h8b: sine = 16'heeef ;
			8'h8c: sine = 16'hed6d ;
			8'h8d: sine = 16'hebed ;
			8'h8e: sine = 16'hea71 ;
			8'h8f: sine = 16'he8f8 ;
			8'h90: sine = 16'he783 ;
			8'h91: sine = 16'he611 ;
			8'h92: sine = 16'he4a4 ;
			8'h93: sine = 16'he33b ;
			8'h94: sine = 16'he1d6 ;
			8'h95: sine = 16'he075 ;
			8'h96: sine = 16'hdf1a ;
			8'h97: sine = 16'hddc4 ;
			8'h98: sine = 16'hdc73 ;
			8'h99: sine = 16'hdb27 ;
			8'h9a: sine = 16'hd9e1 ;
			8'h9b: sine = 16'hd8a1 ;
			8'h9c: sine = 16'hd767 ;
			8'h9d: sine = 16'hd634 ;
			8'h9e: sine = 16'hd506 ;
			8'h9f: sine = 16'hd3e0 ;
			8'ha0: sine = 16'hd2c0 ;
			8'ha1: sine = 16'hd1a7 ;
			8'ha2: sine = 16'hd095 ;
			8'ha3: sine = 16'hcf8b ;
			8'ha4: sine = 16'hce88 ;
			8'ha5: sine = 16'hcd8d ;
			8'ha6: sine = 16'hcc9a ;
			8'ha7: sine = 16'hcbae ;
			8'ha8: sine = 16'hcacb ;
			8'ha9: sine = 16'hc9ef ;
			8'haa: sine = 16'hc91c ;
			8'hab: sine = 16'hc852 ;
			8'hac: sine = 16'hc790 ;
			8'had: sine = 16'hc6d7 ;
			8'hae: sine = 16'hc626 ;
			8'haf: sine = 16'hc57f ;
			8'hb0: sine = 16'hc4e1 ;
			8'hb1: sine = 16'hc44b ;
			8'hb2: sine = 16'hc3bf ;
			8'hb3: sine = 16'hc33c ;
			8'hb4: sine = 16'hc2c3 ;
			8'hb5: sine = 16'hc253 ;
			8'hb6: sine = 16'hc1ec ;
			8'hb7: sine = 16'hc190 ;
			8'hb8: sine = 16'hc13c ;
			8'hb9: sine = 16'hc0f3 ;
			8'hba: sine = 16'hc0b3 ;
			8'hbb: sine = 16'hc07d ;
			8'hbc: sine = 16'hc050 ;
			8'hbd: sine = 16'hc02e ;
			8'hbe: sine = 16'hc015 ;
			8'hbf: sine = 16'hc006 ;
			8'hc0: sine = 16'hc001 ;
			8'hc1: sine = 16'hc006 ;
			8'hc2: sine = 16'hc015 ;
			8'hc3: sine = 16'hc02e ;
			8'hc4: sine = 16'hc050 ;
			8'hc5: sine = 16'hc07d ;
			8'hc6: sine = 16'hc0b3 ;
			8'hc7: sine = 16'hc0f3 ;
			8'hc8: sine = 16'hc13c ;
			8'hc9: sine = 16'hc190 ;
			8'hca: sine = 16'hc1ec ;
			8'hcb: sine = 16'hc253 ;
			8'hcc: sine = 16'hc2c3 ;
			8'hcd: sine = 16'hc33c ;
			8'hce: sine = 16'hc3bf ;
			8'hcf: sine = 16'hc44b ;
			8'hd0: sine = 16'hc4e1 ;
			8'hd1: sine = 16'hc57f ;
			8'hd2: sine = 16'hc626 ;
			8'hd3: sine = 16'hc6d7 ;
			8'hd4: sine = 16'hc790 ;
			8'hd5: sine = 16'hc852 ;
			8'hd6: sine = 16'hc91c ;
			8'hd7: sine = 16'hc9ef ;
			8'hd8: sine = 16'hcacb ;
			8'hd9: sine = 16'hcbae ;
			8'hda: sine = 16'hcc9a ;
			8'hdb: sine = 16'hcd8d ;
			8'hdc: sine = 16'hce88 ;
			8'hdd: sine = 16'hcf8b ;
			8'hde: sine = 16'hd095 ;
			8'hdf: sine = 16'hd1a7 ;
			8'he0: sine = 16'hd2c0 ;
			8'he1: sine = 16'hd3e0 ;
			8'he2: sine = 16'hd506 ;
			8'he3: sine = 16'hd634 ;
			8'he4: sine = 16'hd767 ;
			8'he5: sine = 16'hd8a1 ;
			8'he6: sine = 16'hd9e1 ;
			8'he7: sine = 16'hdb27 ;
			8'he8: sine = 16'hdc73 ;
			8'he9: sine = 16'hddc4 ;
			8'hea: sine = 16'hdf1a ;
			8'heb: sine = 16'he075 ;
			8'hec: sine = 16'he1d6 ;
			8'hed: sine = 16'he33b ;
			8'hee: sine = 16'he4a4 ;
			8'hef: sine = 16'he611 ;
			8'hf0: sine = 16'he783 ;
			8'hf1: sine = 16'he8f8 ;
			8'hf2: sine = 16'hea71 ;
			8'hf3: sine = 16'hebed ;
			8'hf4: sine = 16'hed6d ;
			8'hf5: sine = 16'heeef ;
			8'hf6: sine = 16'hf074 ;
			8'hf7: sine = 16'hf1fb ;
			8'hf8: sine = 16'hf384 ;
			8'hf9: sine = 16'hf510 ;
			8'hfa: sine = 16'hf69d ;
			8'hfb: sine = 16'hf82b ;
			8'hfc: sine = 16'hf9bb ;
			8'hfd: sine = 16'hfb4b ;
			8'hfe: sine = 16'hfcdd ;
			8'hff: sine = 16'hfe6e ;
	endcase
end
endmodule