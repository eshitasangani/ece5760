

module DE1_SoC_Computer (
	////////////////////////////////////
	// FPGA Pins
	////////////////////////////////////

	// Clock pins
	CLOCK_50,
	CLOCK2_50,
	CLOCK3_50,
	CLOCK4_50,

	// ADC
	ADC_CS_N,
	ADC_DIN,
	ADC_DOUT,
	ADC_SCLK,

	// Audio
	AUD_ADCDAT,
	AUD_ADCLRCK,
	AUD_BCLK,
	AUD_DACDAT,
	AUD_DACLRCK,
	AUD_XCK,

	// SDRAM
	DRAM_ADDR,
	DRAM_BA,
	DRAM_CAS_N,
	DRAM_CKE,
	DRAM_CLK,
	DRAM_CS_N,
	DRAM_DQ,
	DRAM_LDQM,
	DRAM_RAS_N,
	DRAM_UDQM,
	DRAM_WE_N,

	// I2C Bus for Configuration of the Audio and Video-In Chips
	FPGA_I2C_SCLK,
	FPGA_I2C_SDAT,

	// 40-Pin Headers
	GPIO_0,
	GPIO_1,
	
	// Seven Segment Displays
	HEX0,
	HEX1,
	HEX2,
	HEX3,
	HEX4,
	HEX5,

	// IR
	IRDA_RXD,
	IRDA_TXD,

	// Pushbuttons
	KEY,

	// LEDs
	LEDR,

	// PS2 Ports
	PS2_CLK,
	PS2_DAT,
	
	PS2_CLK2,
	PS2_DAT2,

	// Slider Switches
	SW,

	// Video-In
	TD_CLK27,
	TD_DATA,
	TD_HS,
	TD_RESET_N,
	TD_VS,

	// VGA
	VGA_B,
	VGA_BLANK_N,
	VGA_CLK,
	VGA_G,
	VGA_HS,
	VGA_R,
	VGA_SYNC_N,
	VGA_VS,

	////////////////////////////////////
	// HPS Pins
	////////////////////////////////////
	
	// DDR3 SDRAM
	HPS_DDR3_ADDR,
	HPS_DDR3_BA,
	HPS_DDR3_CAS_N,
	HPS_DDR3_CKE,
	HPS_DDR3_CK_N,
	HPS_DDR3_CK_P,
	HPS_DDR3_CS_N,
	HPS_DDR3_DM,
	HPS_DDR3_DQ,
	HPS_DDR3_DQS_N,
	HPS_DDR3_DQS_P,
	HPS_DDR3_ODT,
	HPS_DDR3_RAS_N,
	HPS_DDR3_RESET_N,
	HPS_DDR3_RZQ,
	HPS_DDR3_WE_N,

	// Ethernet
	HPS_ENET_GTX_CLK,
	HPS_ENET_INT_N,
	HPS_ENET_MDC,
	HPS_ENET_MDIO,
	HPS_ENET_RX_CLK,
	HPS_ENET_RX_DATA,
	HPS_ENET_RX_DV,
	HPS_ENET_TX_DATA,
	HPS_ENET_TX_EN,

	// Flash
	HPS_FLASH_DATA,
	HPS_FLASH_DCLK,
	HPS_FLASH_NCSO,

	// Accelerometer
	HPS_GSENSOR_INT,
		
	// General Purpose I/O
	HPS_GPIO,
		
	// I2C
	HPS_I2C_CONTROL,
	HPS_I2C1_SCLK,
	HPS_I2C1_SDAT,
	HPS_I2C2_SCLK,
	HPS_I2C2_SDAT,

	// Pushbutton
	HPS_KEY,

	// LED
	HPS_LED,
		
	// SD Card
	HPS_SD_CLK,
	HPS_SD_CMD,
	HPS_SD_DATA,

	// SPI
	HPS_SPIM_CLK,
	HPS_SPIM_MISO,
	HPS_SPIM_MOSI,
	HPS_SPIM_SS,

	// UART
	HPS_UART_RX,
	HPS_UART_TX,

	// USB
	HPS_CONV_USB_N,
	HPS_USB_CLKOUT,
	HPS_USB_DATA,
	HPS_USB_DIR,
	HPS_USB_NXT,
	HPS_USB_STP
);

//=======================================================
//  PARAMETER declarations
//=======================================================


//=======================================================
//  PORT declarations
//=======================================================

////////////////////////////////////
// FPGA Pins
////////////////////////////////////

// Clock pins
input						CLOCK_50;
input						CLOCK2_50;
input						CLOCK3_50;
input						CLOCK4_50;

// ADC
inout						ADC_CS_N;
output					ADC_DIN;
input						ADC_DOUT;
output					ADC_SCLK;

// Audio
input						AUD_ADCDAT;
inout						AUD_ADCLRCK;
inout						AUD_BCLK;
output					AUD_DACDAT;
inout						AUD_DACLRCK;
output					AUD_XCK;

// SDRAM
output 		[12: 0]	DRAM_ADDR;
output		[ 1: 0]	DRAM_BA;
output					DRAM_CAS_N;
output					DRAM_CKE;
output					DRAM_CLK;
output					DRAM_CS_N;
inout			[15: 0]	DRAM_DQ;
output					DRAM_LDQM;
output					DRAM_RAS_N;
output					DRAM_UDQM;
output					DRAM_WE_N;

// I2C Bus for Configuration of the Audio and Video-In Chips
output					FPGA_I2C_SCLK;
inout						FPGA_I2C_SDAT;

// 40-pin headers
inout			[35: 0]	GPIO_0;
inout			[35: 0]	GPIO_1;

// Seven Segment Displays
output		[ 6: 0]	HEX0;
output		[ 6: 0]	HEX1;
output		[ 6: 0]	HEX2;
output		[ 6: 0]	HEX3;
output		[ 6: 0]	HEX4;
output		[ 6: 0]	HEX5;

// IR
input						IRDA_RXD;
output					IRDA_TXD;

// Pushbuttons
input			[ 3: 0]	KEY;

// LEDs
output		[ 9: 0]	LEDR;

// PS2 Ports
inout						PS2_CLK;
inout						PS2_DAT;

inout						PS2_CLK2;
inout						PS2_DAT2;

// Slider Switches
input			[ 9: 0]	SW;

// Video-In
input						TD_CLK27;
input			[ 7: 0]	TD_DATA;
input						TD_HS;
output					TD_RESET_N;
input						TD_VS;

// VGA
output		[ 7: 0]	VGA_B;
output					VGA_BLANK_N;
output					VGA_CLK;
output		[ 7: 0]	VGA_G;
output					VGA_HS;
output		[ 7: 0]	VGA_R;
output					VGA_SYNC_N;
output					VGA_VS;



////////////////////////////////////
// HPS Pins
////////////////////////////////////
	
// DDR3 SDRAM
output		[14: 0]	HPS_DDR3_ADDR;
output		[ 2: 0]  HPS_DDR3_BA;
output					HPS_DDR3_CAS_N;
output					HPS_DDR3_CKE;
output					HPS_DDR3_CK_N;
output					HPS_DDR3_CK_P;
output					HPS_DDR3_CS_N;
output		[ 3: 0]	HPS_DDR3_DM;
inout			[31: 0]	HPS_DDR3_DQ;
inout			[ 3: 0]	HPS_DDR3_DQS_N;
inout			[ 3: 0]	HPS_DDR3_DQS_P;
output					HPS_DDR3_ODT;
output					HPS_DDR3_RAS_N;
output					HPS_DDR3_RESET_N;
input						HPS_DDR3_RZQ;
output					HPS_DDR3_WE_N;

// Ethernet
output					HPS_ENET_GTX_CLK;
inout						HPS_ENET_INT_N;
output					HPS_ENET_MDC;
inout						HPS_ENET_MDIO;
input						HPS_ENET_RX_CLK;
input			[ 3: 0]	HPS_ENET_RX_DATA;
input						HPS_ENET_RX_DV;
output		[ 3: 0]	HPS_ENET_TX_DATA;
output					HPS_ENET_TX_EN;

// Flash
inout			[ 3: 0]	HPS_FLASH_DATA;
output					HPS_FLASH_DCLK;
output					HPS_FLASH_NCSO;

// Accelerometer
inout						HPS_GSENSOR_INT;

// General Purpose I/O
inout			[ 1: 0]	HPS_GPIO;

// I2C
inout						HPS_I2C_CONTROL;
inout						HPS_I2C1_SCLK;
inout						HPS_I2C1_SDAT;
inout						HPS_I2C2_SCLK;
inout						HPS_I2C2_SDAT;

// Pushbutton
inout						HPS_KEY;

// LED
inout						HPS_LED;

// SD Card
output					HPS_SD_CLK;
inout						HPS_SD_CMD;
inout			[ 3: 0]	HPS_SD_DATA;

// SPI
output					HPS_SPIM_CLK;
input						HPS_SPIM_MISO;
output					HPS_SPIM_MOSI;
inout						HPS_SPIM_SS;

// UART
input						HPS_UART_RX;
output					HPS_UART_TX;

// USB
inout						HPS_CONV_USB_N;
input						HPS_USB_CLKOUT;
inout			[ 7: 0]	HPS_USB_DATA;
input						HPS_USB_DIR;
input						HPS_USB_NXT;
output					HPS_USB_STP;

//=======================================================
//  REG/WIRE declarations
//=======================================================

wire			[15: 0]	hex3_hex0;
//wire			[15: 0]	hex5_hex4;

//assign HEX0 = ~hex3_hex0[ 6: 0]; // hex3_hex0[ 6: 0]; 
//assign HEX1 = ~hex3_hex0[14: 8];
//assign HEX2 = ~hex3_hex0[22:16];
//assign HEX3 = ~hex3_hex0[30:24];
assign HEX4 = 7'b1111111;
assign HEX5 = 7'b1111111;

HexDigit Digit0(HEX0, hex3_hex0[3:0]);
HexDigit Digit1(HEX1, hex3_hex0[7:4]);
HexDigit Digit2(HEX2, hex3_hex0[11:8]);
HexDigit Digit3(HEX3, hex3_hex0[15:12]);


//=======================================================
//  DIFFUSION SOLVER
//=======================================================

// PIO //
wire reset_from_hps;
wire pio_done_send;


// m10k //
reg  [18:0] write_addr_u_curr;
reg  [18:0] write_addr_v_next;

reg  [18:0] read_addr_u_curr;
reg  [18:0] read_addr_v_next;

reg         write_en_u_curr;
reg         write_en_v_next;

reg  signed [17:0] write_data_u_curr;
reg  signed [17:0] write_data_v_next;

wire signed [17:0] read_data_u_curr;
wire signed [17:0] read_data_v_next;

// inputs to diffusion solver

reg signed [17:0] v_next;
reg signed [17:0] v_next_reg; // store curr node v_next so we can free solver to calc diffuion of cell above us
reg signed [17:0] u_curr;
reg signed [17:0] u_neighbor_t;
reg signed [17:0] u_neighbor_b;
reg signed [17:0] u_neighbor_l;
reg signed [17:0] u_neighbor_r;
reg signed [17:0] u_neighbor_lc;
reg signed [17:0] u_neighbor_rc;

wire signed [17:0] pio_alpha;
wire signed [17:0] pio_beta;
wire signed [17:0] pio_gamma;

reg  signed [17:0] alpha;
reg  signed [17:0] beta;
reg  signed [17:0] gamma;

// outputs from diffusion solver
wire signed [17:0] u_next_top;
reg  signed [17:0] u_next_reg; // this will store our current node's output so that we can free up the solver to calculate the diffusion of the cell above us. 

wire is_frozen;
reg  is_frozen_reg; // store frozen val for the current node so we can free up solver to calculate diffusion for the node above us.
reg  is_frozen_bottom; // store frozen val for the cell below us 
reg [18:0] is_frozen_y;
reg 	   is_frozen_pio;

/*
neighbor indexing: 
    even:
        4 0 5 
        2 x 3
        - 1 -
    odd:
        - 0 - 
        2 x 3
        4 1 5
*/

diffusion_solver curr_cell (
    .u_neighbor_0 (u_neighbor_t), // top
    .u_neighbor_1 (u_neighbor_b), // bottom
    .u_neighbor_2 (beta),         // left
    .u_neighbor_3 (beta),         // right
    .u_neighbor_4 (beta),         // left corner
    .u_neighbor_5 (beta),         // right corner
    .u_curr       (u_curr),
    .v_next       (v_next),
    .alpha        (alpha),
    .beta         (beta),
      
    .u_next       (u_next_top),
    .is_frozen    (is_frozen)
);

M10K_1000_8 M10k_u_curr ( 
    .q             (read_data_u_curr), 
    .d             (write_data_u_curr), 
    .write_address (write_addr_u_curr),
    .read_address  (read_addr_u_curr),
    .we            (write_en_u_curr),
    .clk           (CLOCK_50)
);

M10K_1000_8 M10k_v_next ( // we only store v_next bc v_next = v_curr + gamma, but we never need to store v_curr
    .q             (read_data_v_next), 
    .d             (write_data_v_next), 
    .write_address (write_addr_v_next),
    .read_address  (read_addr_v_next),
    .we            (write_en_v_next),
    .clk           (CLOCK_50)
);

// ------------------------- //
//       STATE MACHINE       //
// ------------------------- //

// 11 nodes

// reg [15:0] idx;

reg [4:0] state;

always @(posedge CLOCK_50) begin
    if (~KEY[0] || reset_from_hps) begin
        write_data_u_curr <= beta;
        write_data_v_next <= 18'd0;
        write_addr_u_curr <= 19'd0;
        write_addr_v_next <= 19'd0;
        write_en_u_curr <= 1'd1;
        write_en_v_next <= 1'd1;

        read_addr_u_curr <= 19'd0;
        read_addr_v_next <= 19'd0;

		alpha <= pio_alpha;
		beta  <= pio_beta;
		gamma <= pio_gamma;

        state  <= 5'd0;
    end
    else begin
        case (state)

            5'd0: begin // initialization
                // SETTING INITIAL U AND V VALUES //
                // only center node is frozen, set to 1
                if (write_addr_u_curr == 19'd3) begin 
                    // on next cycle, it'll be the center node
                    write_data_u_curr <= 18'd0;
                    write_data_v_next <= 18'b01_0000000000000000 + gamma;
                end
                else if (write_addr_u_curr == 19'd2 || write_addr_u_curr == 19'd4) begin
                    // the nodes around the center node are receptive, but not frozen 
                    write_data_u_curr <= 18'd0;
                    write_data_v_next <= beta + gamma;
                end
                else begin
                    // all other nodes are nonreceptive
                    write_data_u_curr <= beta;
                    write_data_v_next <= 18'd0;
                end

                // MOVE FORWARD OR STOP //
                if (write_addr_u_curr >= 19'd10) begin
                    state <= 5'd1;
                    write_addr_u_curr <= 19'd0;
                    write_addr_v_next <= 19'd0;
                    write_en_u_curr <= 1'd0;
                    write_en_v_next <= 1'd0;
                end
                else begin
                    state <= 5'd0;
                    write_addr_u_curr <= write_addr_u_curr + 19'd1;
                    write_addr_v_next <= write_addr_v_next + 19'd1;
                    write_en_u_curr <= 1'd1;
                    write_en_v_next <= 1'd1;
                end
            end

            5'd1: begin
                u_neighbor_b      <= beta; // bottom 

                // read from m10ks for u_curr and v_next for this cell
                u_curr            <= read_data_u_curr;
                v_next            <= ((read_data_v_next + gamma) >= 18'b01_0000000000000000)? 18'b01_0000000000000000 : (read_data_v_next + gamma);
                read_addr_u_curr  <= read_addr_u_curr + 19'd1;
                state             <= 5'd2;
            end

            5'd2: begin
                // wait for next read to come back
                state             <= 5'd3;
            end
            5'd3: begin
                // read from m10k for top neighbor
                u_neighbor_t <= read_data_u_curr; 

                // increment these now, so we can read them a cycle earlier
                read_addr_u_curr <= read_addr_u_curr + 19'd1;
                read_addr_v_next <= read_addr_v_next + 19'd1;

                state             <= 5'd4;
            end
            5'd4: begin
				if (pio_done_send) begin // we have to wait for the hps to request the next value
					// now we can use diffusion solver output
					// store these outputs and then move up to calculate diffusion for the cell above us. 
					is_frozen_reg <= is_frozen;
					is_frozen_y   <= write_addr_u_curr;
					is_frozen_pio <= is_frozen;

					u_next_reg <= u_next_top; // u_next_top is solver output
					v_next_reg <= v_next;                

					// take a step up
					u_neighbor_b <= u_curr;
					u_curr <= u_neighbor_t;
                	state <= 5'd5;
				end
				else begin
					state <= 5'd4;
				end
            end
            5'd5: begin // read m10k for the cell above us so we can calc diffusion for it
				if (!pio_done_send) begin
					// read from m10k for top neighbor
					u_neighbor_t <= read_data_u_curr; 

					// read from m10k for v_next
					v_next            <= ((read_data_v_next + gamma) >= 18'b01_0000000000000000)? 18'b01_0000000000000000 : (read_data_v_next + gamma);

					// increment these now, so we can read them a cycle earlier
					read_addr_u_curr <= read_addr_u_curr + 19'd1;
					read_addr_v_next <= read_addr_v_next + 19'd1;

					state             <= 5'd6;
				end
				else begin
					state <= 5'd5;
				end

            end
            5'd6: begin
				if (!pio_done_send) begin
					// check if any neighbors are frozen
					// eventually will have to also check r,l,rc,rl neighbors too but 
					// right now r,l,rc,rl are edge cells so they are static
					if (is_frozen_reg || is_frozen_bottom || is_frozen) begin
						// if we or any neighbors are frozen, we are a receptive cell.
						// write the new s=u+v value to v, write 0 to u
						write_data_v_next <= v_next_reg + u_next_reg;
						write_data_u_curr <= 18'd0;
					end
					else begin
						// if us and none of our neighbors are frozen, we are a non-receptive cell
						// write 0 to v, write the new s=u+v value to u
						write_data_v_next <= 18'd0;
						write_data_u_curr <= v_next_reg + u_next_reg;
					end

					write_en_u_curr <= 1'b1;
					write_en_v_next <= 1'b1;

					state <= 5'd7;
				end
				else begin
					state <= 5'd6;
				end
            end
            5'd7: begin
				if (pio_done_send) begin // we have to wait for the hps to request the next value
                	// move up one cell!
					u_neighbor_b <= u_curr;
					u_curr       <= u_neighbor_t;

					is_frozen_bottom <= is_frozen_reg;
					is_frozen_reg    <= is_frozen;
					is_frozen_y      <= write_addr_u_curr + 19'd1;
					is_frozen_pio    <= is_frozen;

					u_next_reg <= u_next_top;
					v_next_reg <= v_next;

					// read from m10k for top neighbor
					u_neighbor_t <= (read_addr_u_curr >= 19'd10) ? beta : read_data_u_curr; // consider top edge boundary

					// read from m10k for v_next
					v_next <= (read_addr_v_next >= 19'd10) ? 18'd0 : (((read_data_v_next + gamma) >= 18'b01_0000000000000000)? 18'b01_0000000000000000 : (read_data_v_next + gamma)); // consider top edge boundary

					// incr write addresses
					if (write_addr_u_curr >= 19'd10) begin
						write_addr_u_curr <= 19'd0;
						write_addr_v_next <= 19'd0;
						read_addr_u_curr  <= 19'd0;
						read_addr_v_next  <= 19'd0;
						state <= 5'd8;
					end
					else begin
						write_addr_u_curr <= write_addr_u_curr + 19'd1;
						write_addr_v_next <= write_addr_v_next + 19'd1;
						// increment these now, so we can read them a cycle earlier
						// consider top edge boundary: make sure we're not trying to read nonexistent data from m10ks
						read_addr_u_curr  <= (read_addr_u_curr >= 19'd10) ? read_addr_u_curr : (read_addr_u_curr + 19'd1);
						read_addr_v_next  <= (read_addr_v_next >= 19'd10) ? read_addr_v_next : (read_addr_v_next + 19'd1);
						state             <= 5'd6;
					end
					write_en_u_curr <= 1'b0;
					write_en_v_next <= 1'b0;
				end
				else begin
					state <= 5'd7;
				end
            end

            5'd8: begin // this is a wait state so we can get our read data at the bottom in state 1 
				if (!pio_done_send) begin
                	state <= 5'd1;
				end
				else begin
					state <= 5'd8;
				end
            end

        endcase
    end
end



//=======================================================
//  Structural coding
//=======================================================

Computer_System The_System (
	////////////////////////////////////
	// FPGA Side
	////////////////////////////////////

	// Global signals
	.system_pll_ref_clk_clk					(CLOCK_50),
	.system_pll_ref_reset_reset			(1'b0),

	// AV Config
	.av_config_SCLK							(FPGA_I2C_SCLK),
	.av_config_SDAT							(FPGA_I2C_SDAT),

	// Slider Switches
	.slider_switches_export					(SW),

	// Pushbuttons (~KEY[3:0]),
	.pushbuttons_export						(~KEY[3:0]),

	// LEDs
	.leds_export								(LEDR),
	
	// Seven Segs
	.hex3_hex0_export							(hex3_hex0),


	// VGA Subsystem
	.vga_pll_ref_clk_clk 					(CLOCK2_50),
	.vga_pll_ref_reset_reset				(1'b0),
	.vga_CLK										(VGA_CLK),
	.vga_BLANK									(VGA_BLANK_N),
	.vga_SYNC									(VGA_SYNC_N),
	.vga_HS										(VGA_HS),
	.vga_VS										(VGA_VS),
	.vga_R										(VGA_R),
	.vga_G										(VGA_G),
	.vga_B										(VGA_B),
	
	
	////////////////////////////////////
	// HPS Side
	////////////////////////////////////
	// DDR3 SDRAM
	.memory_mem_a			(HPS_DDR3_ADDR),
	.memory_mem_ba			(HPS_DDR3_BA),
	.memory_mem_ck			(HPS_DDR3_CK_P),
	.memory_mem_ck_n		(HPS_DDR3_CK_N),
	.memory_mem_cke		(HPS_DDR3_CKE),
	.memory_mem_cs_n		(HPS_DDR3_CS_N),
	.memory_mem_ras_n		(HPS_DDR3_RAS_N),
	.memory_mem_cas_n		(HPS_DDR3_CAS_N),
	.memory_mem_we_n		(HPS_DDR3_WE_N),
	.memory_mem_reset_n	(HPS_DDR3_RESET_N),
	.memory_mem_dq			(HPS_DDR3_DQ),
	.memory_mem_dqs		(HPS_DDR3_DQS_P),
	.memory_mem_dqs_n		(HPS_DDR3_DQS_N),
	.memory_mem_odt		(HPS_DDR3_ODT),
	.memory_mem_dm			(HPS_DDR3_DM),
	.memory_oct_rzqin		(HPS_DDR3_RZQ),
		  
	// Ethernet
	.hps_io_hps_io_gpio_inst_GPIO35	(HPS_ENET_INT_N),
	.hps_io_hps_io_emac1_inst_TX_CLK	(HPS_ENET_GTX_CLK),
	.hps_io_hps_io_emac1_inst_TXD0	(HPS_ENET_TX_DATA[0]),
	.hps_io_hps_io_emac1_inst_TXD1	(HPS_ENET_TX_DATA[1]),
	.hps_io_hps_io_emac1_inst_TXD2	(HPS_ENET_TX_DATA[2]),
	.hps_io_hps_io_emac1_inst_TXD3	(HPS_ENET_TX_DATA[3]),
	.hps_io_hps_io_emac1_inst_RXD0	(HPS_ENET_RX_DATA[0]),
	.hps_io_hps_io_emac1_inst_MDIO	(HPS_ENET_MDIO),
	.hps_io_hps_io_emac1_inst_MDC		(HPS_ENET_MDC),
	.hps_io_hps_io_emac1_inst_RX_CTL	(HPS_ENET_RX_DV),
	.hps_io_hps_io_emac1_inst_TX_CTL	(HPS_ENET_TX_EN),
	.hps_io_hps_io_emac1_inst_RX_CLK	(HPS_ENET_RX_CLK),
	.hps_io_hps_io_emac1_inst_RXD1	(HPS_ENET_RX_DATA[1]),
	.hps_io_hps_io_emac1_inst_RXD2	(HPS_ENET_RX_DATA[2]),
	.hps_io_hps_io_emac1_inst_RXD3	(HPS_ENET_RX_DATA[3]),

	// Flash
	.hps_io_hps_io_qspi_inst_IO0	(HPS_FLASH_DATA[0]),
	.hps_io_hps_io_qspi_inst_IO1	(HPS_FLASH_DATA[1]),
	.hps_io_hps_io_qspi_inst_IO2	(HPS_FLASH_DATA[2]),
	.hps_io_hps_io_qspi_inst_IO3	(HPS_FLASH_DATA[3]),
	.hps_io_hps_io_qspi_inst_SS0	(HPS_FLASH_NCSO),
	.hps_io_hps_io_qspi_inst_CLK	(HPS_FLASH_DCLK),

	// Accelerometer
	.hps_io_hps_io_gpio_inst_GPIO61	(HPS_GSENSOR_INT),


	// General Purpose I/O
	.hps_io_hps_io_gpio_inst_GPIO40	(HPS_GPIO[0]),
	.hps_io_hps_io_gpio_inst_GPIO41	(HPS_GPIO[1]),

	// I2C
	.hps_io_hps_io_gpio_inst_GPIO48	(HPS_I2C_CONTROL),
	.hps_io_hps_io_i2c0_inst_SDA		(HPS_I2C1_SDAT),
	.hps_io_hps_io_i2c0_inst_SCL		(HPS_I2C1_SCLK),
	.hps_io_hps_io_i2c1_inst_SDA		(HPS_I2C2_SDAT),
	.hps_io_hps_io_i2c1_inst_SCL		(HPS_I2C2_SCLK),

	// Pushbutton
	.hps_io_hps_io_gpio_inst_GPIO54	(HPS_KEY),

	// LED
	.hps_io_hps_io_gpio_inst_GPIO53	(HPS_LED),

	// SD Card
	.hps_io_hps_io_sdio_inst_CMD	(HPS_SD_CMD),
	.hps_io_hps_io_sdio_inst_D0	(HPS_SD_DATA[0]),
	.hps_io_hps_io_sdio_inst_D1	(HPS_SD_DATA[1]),
	.hps_io_hps_io_sdio_inst_CLK	(HPS_SD_CLK),
	.hps_io_hps_io_sdio_inst_D2	(HPS_SD_DATA[2]),
	.hps_io_hps_io_sdio_inst_D3	(HPS_SD_DATA[3]),

	// SPI
	.hps_io_hps_io_spim1_inst_CLK		(HPS_SPIM_CLK),
	.hps_io_hps_io_spim1_inst_MOSI	(HPS_SPIM_MOSI),
	.hps_io_hps_io_spim1_inst_MISO	(HPS_SPIM_MISO),
	.hps_io_hps_io_spim1_inst_SS0		(HPS_SPIM_SS),

	// UART
	.hps_io_hps_io_uart0_inst_RX	(HPS_UART_RX),
	.hps_io_hps_io_uart0_inst_TX	(HPS_UART_TX),

	// USB
	.hps_io_hps_io_gpio_inst_GPIO09	(HPS_CONV_USB_N),
	.hps_io_hps_io_usb1_inst_D0		(HPS_USB_DATA[0]),
	.hps_io_hps_io_usb1_inst_D1		(HPS_USB_DATA[1]),
	.hps_io_hps_io_usb1_inst_D2		(HPS_USB_DATA[2]),
	.hps_io_hps_io_usb1_inst_D3		(HPS_USB_DATA[3]),
	.hps_io_hps_io_usb1_inst_D4		(HPS_USB_DATA[4]),
	.hps_io_hps_io_usb1_inst_D5		(HPS_USB_DATA[5]),
	.hps_io_hps_io_usb1_inst_D6		(HPS_USB_DATA[6]),
	.hps_io_hps_io_usb1_inst_D7		(HPS_USB_DATA[7]),
	.hps_io_hps_io_usb1_inst_CLK		(HPS_USB_CLKOUT),
	.hps_io_hps_io_usb1_inst_STP		(HPS_USB_STP),
	.hps_io_hps_io_usb1_inst_DIR		(HPS_USB_DIR),
	.hps_io_hps_io_usb1_inst_NXT		(HPS_USB_NXT),

	// PIO
	.pio_done_send_external_connection_export      (pio_done_send),
	.pio_reset_to_hps_external_connection_export   (~KEY[0]),   //   pio_reset_to_hps_external_connection.export
	.pio_reset_from_hps_external_connection_export (reset_from_hps), // pio_reset_from_hps_external_connection.export
	.is_frozen_y_external_connection_export        (is_frozen_y),        //        is_frozen_y_external_connection.export
	.is_frozen_pio_external_connection_export      (is_frozen_pio),        //        is_frozen_x_external_connection.export
	.pio_gamma_external_connection_export          (pio_gamma),          //          pio_gamma_external_connection.export
	.pio_beta_external_connection_export           (pio_beta),           //           pio_beta_external_connection.export
	.pio_alpha_external_connection_export          (pio_alpha)           //          pio_alpha_external_connection.export
);

endmodule

/*
    this module calculates the diffusion equation (u) of one cell 
    it also outputs whether this cell is frozen at the end of calculating the diffusion
    u_next = u_curr + alpha / 2 * (u_avg - u_curr)
    u_avg = avg u over all neighbors
*/
module diffusion_solver (
    input  wire signed [17:0] u_neighbor_0,
    input  wire signed [17:0] u_neighbor_1,
    input  wire signed [17:0] u_neighbor_2,
    input  wire signed [17:0] u_neighbor_3,
    input  wire signed [17:0] u_neighbor_4,
    input  wire signed [17:0] u_neighbor_5,
    input  wire signed [17:0] u_curr,
    input  wire signed [17:0] v_next, // this is calculated outside of this module, when we calculate our current u and v

    input  wire signed [17:0] alpha,
    input  wire signed [17:0] beta,

    output wire signed [17:0] u_next,

    output wire        is_frozen
);

    wire signed [17:0] u_avg_0;
    wire signed [17:0] u_avg_1;
    wire signed [17:0] u_avg_total;
    wire signed [17:0] laplace_out;
    wire signed [17:0] u_next_tmp;

    // s = u + v
    // frozen if s >= 1
    assign is_frozen = ((u_next + v_next) >= 18'b01_0000000000000000);
    assign u_next_tmp = (u_curr + laplace_out); 
    assign u_next = (u_next_tmp >= 18'b01_0000000000000000) ? 18'b01_0000000000000000 : u_next_tmp;

    signed_mult u_avg_calc0 ( // divide by 6 (num neighbors) -- mult by 1/6
        .out(u_avg_0),
        .a  (u_neighbor_0+u_neighbor_1+u_neighbor_2),
        .b  (18'b00_0010101010101010) // 1/6
    );

    signed_mult u_avg_calc1 ( // divide by 6 (num neighbors) -- mult by 1/6
        .out(u_avg_1),
        .a  (u_neighbor_3+u_neighbor_4+u_neighbor_5),
        .b  (18'b00_0010101010101010) // 1/6
    );

    assign u_avg_total = u_avg_0 + u_avg_1;

    signed_mult laplace_calc ( // alpha / 2 * (u_avg - cell.u)
        .out(laplace_out),
        .a  (alpha >>> 1),
        .b  (u_avg_total - u_curr)
    );

endmodule

//////////////////////////////////////////////////
//// signed mult of 2.16 format 2'comp////////////
//////////////////////////////////////////////////

module signed_mult (out, a, b);
	output 	signed  [17:0]	out;
	input 	signed	[17:0] 	a;
	input 	signed	[17:0] 	b;
	// intermediate full bit length
	wire 	signed	[35:0]	mult_out;
	assign mult_out = a * b;
	// select bits for 7.20 fixed point
	assign out = {mult_out[35], mult_out[34:16]};
endmodule
//////////////////////////////////////////////////


//============================================================
// M10K module for testing
//============================================================
// See example 12-16 in 
// http://people.ece.cornell.edu/land/courses/ece5760/DE1_SOC/HDL_style_qts_qii51007.pdf
//============================================================

module M10K_1000_8( 
    output reg [17:0] q,
    input [17:0] d,
    input [18:0] write_address, read_address,
    input we, clk
);
	 // force M10K ram style
    reg [17:0] mem [10:0]  /* synthesis ramstyle = "no_rw_check, M10K" */;
    always @ (posedge clk) begin
        if (we) begin
            mem[write_address] <= d;
		  end
        q <= mem[read_address]; // q doesn't get d in this clock cycle
    end
endmodule